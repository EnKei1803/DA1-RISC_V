module CONTROL_UNIT
#(parameter n = 32)
(
	input [n-1:0] Din,
	
input  clk,
input  [8:0] IRin,
input  [0:0] run, rstn,
output  [7:0] sel_out, 	//R0->R7 out
output  [0:0] Gout,DINout, //out
output  [0:0] done,
output  [7:0] sel_in, 
output  [0:0] Ain, addsub,Gin,	//R0->7  in
output  [0:0] IRin_en
);



/*

// Control FSM flip-flops 
always_ff @ ( posedge clk , negedge rstn ) begin
if ( !rstn )
state_reg <= T0 ;
else
state_reg <= state_next ;
end

// state register
typedef enum logic[1:0] {T0 = 2'b00, T1 = 2'b01, T2 = 2'b10, T3 = 2'b11} states ; 
states state_reg;
states state_next;

// Control FSM state table 
always_comb begin 
	case (state_reg) 
	T0:
		if (!run & done) state_next = T0; 
		else state_next = T1; 

	T1: 
		if (done) state_next = T0; 
		else state_next = T2; 

	T2:
		state_next = T3; 

	T3: 
		state_next = T0; 
	endcase 
end 



// Control FSM outputs 
	//Choose function
	
logic 	[3:0] temp4;

assign I = IRin[8:6]; 

localparam mv  = 3'b000;	// Rx <- [Ry]
localparam mvi = 3'b001;	// Rx <- DIN[2:0]   
localparam add = 3'b010;	// Rx <- [Rx] + [Ry]
localparam sub = 3'b011;	// Rx <- [Rx] - [Ry]

*/









endmodule
















