
//--------------------------------SHIFTER_32bits------------------------------------
/*
			|--------------------|-----------|-----------|-----------|
			|	 OPERATING MODE	|		S2		|		s1		|		S0		|
			|--------------------|-----------|-----------|-----------|
			|			LOCKED		|		0		|		0		|		0		|
			|--------------------|-----------|-----------|-----------|
			|		SHIFT RIGHT		|		0		|		1		|		0		|
			|--------------------|-----------|-----------|-----------|
			|		SHIFT LEFT		|		1		|		0		|		0		|
			|--------------------|-----------|-----------|-----------|
			|	PARALLEL LOADING	|		1		|		1		|		0		|
			|--------------------|-----------|-----------|-----------|
			|			 ASR			|		0		|		0		|		1		|
			|--------------------|-----------|-----------|-----------|
			|			 ASL			|		0		|		1		|		1		|
			|--------------------|-----------|-----------|-----------|
			|		Rotate Right	|		1		|		0		|		1		|
			|--------------------|-----------|-----------|-----------|
			|		Rotate Left		|		1		|		1		|		1		|
			|--------------------|-----------|-----------|-----------|

*/
module UNIVERSAL_SHIFTER
#(parameter n = 32)
(
	input [n-1:0] 	I,
	input [1:0] 	S,
	input clk, resetn,
	output reg [n-1:0] A
);
	
logic [n-1:0] B;
logic ze_0, ze_1;
assign ze_0 = 1'b0;
assign ze_1 = 1'b0;

REG_32bits_noEN REG_32bits_noEN_1 (B, clk, resetn, A);

//							S1 S0    I0      I1     I2     I3     Y
MUX_4x1 MUX_4x1_01 (S[1:0],  A[0],  A[1],  ze_0,  I[0],  B[0]);
MUX_4x1 MUX_4x1_02 (S[1:0],  A[1],  A[2],  A[0],  I[1],  B[1]);
MUX_4x1 MUX_4x1_03 (S[1:0],  A[2],  A[3],  A[1],  I[2],  B[2]);
MUX_4x1 MUX_4x1_04 (S[1:0],  A[3],  A[4],  A[2],  I[3],  B[3]);
MUX_4x1 MUX_4x1_05 (S[1:0],  A[4],  A[5],  A[3],  I[4],  B[4]);
MUX_4x1 MUX_4x1_06 (S[1:0],  A[5],  A[6],  A[4],  I[5],  B[5]);
MUX_4x1 MUX_4x1_07 (S[1:0],  A[6],  A[7],  A[5],  I[6],  B[6]);
MUX_4x1 MUX_4x1_08 (S[1:0],  A[7],  A[8],  A[6],  I[7],  B[7]);
 
MUX_4x1 MUX_4x1_09 (S[1:0],  A[8],  A[9],  A[7],  I[8],  B[8]);
MUX_4x1 MUX_4x1_10 (S[1:0],  A[9], A[10],  A[8],  I[9],  B[9]);
MUX_4x1 MUX_4x1_11 (S[1:0], A[10], A[11],  A[9], I[10], B[10]);
MUX_4x1 MUX_4x1_12 (S[1:0], A[11], A[12], A[10], I[11], B[11]);
MUX_4x1 MUX_4x1_13 (S[1:0], A[12], A[13], A[11], I[12], B[12]);
MUX_4x1 MUX_4x1_14 (S[1:0], A[13], A[14], A[12], I[13], B[13]);
MUX_4x1 MUX_4x1_15 (S[1:0], A[14], A[15], A[13], I[14], B[14]);
MUX_4x1 MUX_4x1_16 (S[1:0], A[15], A[16], A[14], I[15], B[15]);

MUX_4x1 MUX_4x1_17 (S[1:0], A[16], A[17], A[15], I[16], B[16]);
MUX_4x1 MUX_4x1_18 (S[1:0], A[17], A[18], A[16], I[17], B[17]);
MUX_4x1 MUX_4x1_19 (S[1:0], A[18], A[19], A[17], I[18], B[18]);
MUX_4x1 MUX_4x1_20 (S[1:0], A[19], A[20], A[18], I[19], B[19]);
MUX_4x1 MUX_4x1_21 (S[1:0], A[20], A[21], A[19], I[20], B[20]);
MUX_4x1 MUX_4x1_22 (S[1:0], A[21], A[22], A[20], I[21], B[21]);
MUX_4x1 MUX_4x1_23 (S[1:0], A[22], A[23], A[21], I[22], B[22]);
MUX_4x1 MUX_4x1_24 (S[1:0], A[23], A[24], A[22], I[23], B[23]);

MUX_4x1 MUX_4x1_25 (S[1:0], A[24], A[25], A[23], I[24], B[24]);
MUX_4x1 MUX_4x1_26 (S[1:0], A[25], A[26], A[24], I[25], B[25]);
MUX_4x1 MUX_4x1_27 (S[1:0], A[26], A[27], A[25], I[26], B[26]);
MUX_4x1 MUX_4x1_28 (S[1:0], A[27], A[28], A[26], I[27], B[27]);
MUX_4x1 MUX_4x1_29 (S[1:0], A[28], A[29], A[27], I[28], B[28]);
MUX_4x1 MUX_4x1_30 (S[1:0], A[29], A[30], A[28], I[29], B[29]);
MUX_4x1 MUX_4x1_31 (S[1:0], A[30], A[31], A[29], I[30], B[30]);
MUX_4x1 MUX_4x1_32 (S[1:0], A[31],  ze_1, A[30], I[31], B[31]);

endmodule 

//--------------------------------MUX 4x1------------------------------------

module MUX_4x1
(
	input [1:0] s,
	input I0, I1, I2, I3,
	output Y
);

assign Y =	 s[1] &  s[0] & I3 |			// [1:0]s = 11			Parallel Loading 
				 s[1] & ~s[0] & I2 |			// [1:0]s = 10			Shift Left
				~s[1] &  s[0] & I1 |			// [1:0]s = 01			Shift Right
				~s[1] & ~s[0] & I0 ;			// [1:0]s = 00			Locked
				
endmodule

//--------------------------------REGISTER without ENABLE------------------------------------

module REG_32bits_noEN 
#(parameter n = 32)
(
	input [n-1:0] R,
	input clk, resetn,
	output reg [n-1:0] Q
);

always @(posedge clk or negedge resetn) begin
	if (!resetn) 						// resetn = 0, REG = 0x00
		Q <= {n{1'b0}};
	else 
		Q <= R;										
end

endmodule
