module BRANCH_COMPARE
(
	input 


);